module seg7nmbr(seg_in,seg_out);
  input [3:0]seg_in;
  output [6:0]seg_out;
   reg [6:0]seg_out;
  always @(seg_in)
    begin
      case(seg_in)
          4'b0000:
            begin 
              seg_out=7'b1000000;
            end
          4'b0001:
            begin 
              seg_out=7'b1111001;
            end
          4'b0010: 
            begin
              seg_out=7'b0100100;
            end
          4'b0011: 
            begin
              seg_out=7'b0110000;
            end
          4'b0100: 
            begin
              seg_out=7'b0011011;
            end
          4'b0101:
            begin 
              seg_out=7'b0010010;
            end
          4'b0110: 
            begin
              seg_out=7'b0000010;
            end
          4'b0111: 
            begin
              seg_out=7'b1111000;
            end
          4'b1000: 
            begin
              seg_out=7'b0000000;
            end
          4'b1001: 
            begin
              seg_out=7'b0011000;
            end
          4'b1010: 
            begin
              seg_out=7'b0001000;
            end
          4'b1011: 
            begin
              seg_out=7'b0000011;
            end
          4'b1100: 
            begin
              seg_out=7'b1000110;
            end
          4'b1101: 
            begin
              seg_out=7'b1000000;
            end
          4'b1110: 
            begin
              seg_out=7'b0000110;
            end
          4'b1111: 
            begin
              seg_out=7'b0001110;
            end
          default:
            begin
              seg_out=7'b1111111;
            end
      endcase
    end
endmodule 
