
module gamecontroller(clk, rst, mode, update, timeout2sec, rain, reqlfsr, req2sec, allowgt, raout1, raout2, raout3, raout4, raout5, segen);
input clk, rst, mode, update, timeout2sec;
input [3:0]rain;
output reg reqlfsr, req2sec, allowgt, segen;
output reg [3:0]raout1, raout2, raout3, raout4, raout5;
parameter init=0, start=1, request1=2, waitc1=4, load1=3, request2=5, waitc2=7, load2=6, request3=8, waitc3=10, load3=9, request4=11, waitc4=13, 
load4=12, request5=14, waitc5=16, load5=15, stop=17;
reg [4:0]state;
always @(posedge clk)
  begin
    if(rst==0)
      begin
        state<=init;
      end
    else
      begin
        case(state)
          init:
            begin
              reqlfsr<=0;
              req2sec<=0;
              allowgt<=0;
              segen<=0;
              raout1<=4'h0;
              raout2<=4'h0;
              raout3<=4'h0;
              raout4<=4'h0;
              raout5<=4'h0;
              if(mode==1)
                begin
                  state<=start;
                end
              else
                begin
                  state<=init;
                end
            end
          start:
            begin
              if(update==1)
                begin
                  allowgt<=0;
                  state<=request1;
                end
              else
                begin
                  state<=start;
                end
            end
          request1:
            begin
              reqlfsr=1'b1;
              segen<=1;
              req2sec<=1;
              state<=load1;
            end
          load1:
            begin
              reqlfsr<=1'b0;
              state<=waitc1;
            end
          waitc1:
            begin
              reqlfsr<=1'b0;
              raout1<=rain;
              if(timeout2sec==1)
                begin
                  req2sec<=0;
                  state<=request2;
                end
              else
                begin
                  state<=waitc1;
                end
            end
          request2:
            begin
              reqlfsr=1'b1;
              segen<=1;
              req2sec<=1;
              state<=load2;
            end
         load2:
            begin
              reqlfsr<=1'b0;
              state<=waitc2;
            end
          waitc2:
            begin
              reqlfsr<=1'b0;
              raout2<=rain;
              if(timeout2sec==1)
                begin
                  req2sec<=0;
                  state<=request3;
                end
              else
                begin
                  state<=waitc2;
                end
            end
          request3:
            begin
              reqlfsr=1'b1;
              segen<=1;
              req2sec<=1;
              state<=load3;
            end
         load3:
            begin
              reqlfsr<=1'b0;
              state<=waitc3;
            end
          waitc3:
            begin
              reqlfsr<=1'b0;
              raout3<=rain;
              if(timeout2sec==1)
                begin
                  req2sec<=0;
                  state<=request4;
                end
              else
                begin
                  state<=waitc3;
                end
            end
          request4:
            begin
              reqlfsr=1'b1;
              segen<=1;
              req2sec<=1;
              state<=load4;
            end
          load4:
            begin
              reqlfsr<=1'b0;
              state<=waitc4;
            end
          waitc4:
            begin
              reqlfsr<=1'b0;
              raout4<=rain;
              if(timeout2sec==1)
                begin
                  req2sec<=0;
                  state<=request5;
                end
              else
                begin
                  state<=waitc4;
                end
            end
          request5:
            begin
              reqlfsr=1'b1;
              segen<=1;
              req2sec<=1;
              state<=load5;
            end
          load5:
            begin
              reqlfsr<=1'b0;
              state<=waitc5;
            end
          waitc5:
            begin
              reqlfsr<=1'b0;
              raout5<=rain;
              if(timeout2sec==1)
                begin
                  req2sec<=0;
                  state<=stop;
                end
              else
                begin
                  state<=waitc5;
                end
            end
          stop:
            begin
              allowgt<=1;
              segen<=0;
              state<=start;
            end
          default:
            begin
              state<=init;
            end
        endcase
      end
  end
endmodule            
              


