module accessctrl(clk, rst, valid, alph1, alph2, alph3, alph4, alph5, playeralph, allow, segen);
input clk, valid, rst;
input [3:0]alph1, alph2, alph3, alph4, alph5, playeralph;
output reg allow, segen;
reg flag_red;
parameter init=0, bit1=1, bit2=2, bit3=3, bit4=4, verify=5;
reg [2:0]state;
  always @(posedge clk)
    begin
      if(rst==0)
        begin
          segen<=0;
          state<=init;
        end
      else
        begin
          case(state)
            init:
              begin
                allow<=1'b0;
                flag_red<=1'b0;
                if(valid==1)
                  begin
                    segen<=1;
                    if(alph1!=playeralph)
                      begin
                        flag_red<=1'b1;
                      end
                    state<=bit1;
                  end
                else
                  begin
                    state<=init;
                  end
              end
            bit1:
              begin
                allow<=1'b0;
                if(valid==1)
                  begin
                    if(alph2!=playeralph)
                      begin
                        flag_red<=1'b1;
                      end
                    state<=bit2;
                  end
                else
                  begin
                    state<=bit1;
                  end
              end
            bit2:
              begin
                allow<=1'b0;
                if(valid==1)
                  begin
                    if(alph3!=playeralph)
                      begin
                        flag_red<=1'b1;
                      end
                    state<=bit3;
                  end
                else
                  begin
                    state<=bit2;
                  end
              end
            bit3:
              begin
                allow<=1'b0;
                if(valid==1)
                  begin
                    if(alph4!=playeralph)
                      begin
                        flag_red<=1'b1;
                      end
                    state<=bit4;
                  end
                else
                  begin
                    state<=bit3;
                  end
              end
            bit4:
              begin
                allow<=1'b0;
                if(valid==1)
                  begin
                    if(alph5!=playeralph)
                      begin
                        flag_red<=1'b1;
                      end
                    state<=verify;
                  end
                else
                  begin
                    state<=bit4;
                  end
              end
            verify:
              begin
                if(flag_red==0)
                  begin
                    allow<=1'b1;
                  end
                else
                  begin
                    allow<=1'b0;
                  end
                state<=init;
              end
            default:
              begin
                allow<=1'b0;
                state<=init;
              end
          endcase
        end
    end
endmodule                                    

 